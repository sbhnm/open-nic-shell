`define KEEP  (* keep="TRUE" *)
`define DEBUG (* mark_debug = "true" *)

