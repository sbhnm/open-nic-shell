`include "pcie_spmv_macros.vh"
`timescale 1ns/1ps

module hbm_ctrl #(
    
) (
    input [32*1-1:0]    AXI_ACLK,
    input [32*1-1:0]    AXI_ARESET_N,
    input [32*33 -1: 0]     AXI_ARADDR,
    input [32*2 -1: 0]      AXI_ARBURST,
    input [32*6 -1: 0]      AXI_ARID,
    input [32*4 -1: 0]      AXI_ARLEN,
    input [32*3 -1: 0]      AXI_ARSIZE,
    input [32*1-1:0]    AXI_ARVALID,
    input [32*33 -1: 0]     AXI_AWADDR,
    input [32*2 -1: 0]      AXI_AWBURST,
    input [32*6 -1: 0]      AXI_AWID,
    input [32*4 -1: 0]      AXI_AWLEN,
    input [32*3 -1: 0]      AXI_AWSIZE,
    input [32*1-1:0]    AXI_AWVALID,
    input [32*1-1:0]    AXI_RREADY,
    input [32*1-1:0]    AXI_BREADY,
    input [32*256 -1: 0]    AXI_WDATA,
    input [32*1-1:0]    AXI_WLAST,
    input [32*32 -1: 0]     AXI_WSTRB,
    input [32*32 -1: 0]     AXI_WDATA_PARITY,
    input [32*1-1:0]    AXI_WVALID,
    output [32*1-1:0]   AXI_ARREADY,
    output [32*1-1:0]   AXI_AWREADY,
    output [32*32 -1: 0]    AXI_RDATA_PARITY,
    output [32*256 -1: 0]   AXI_RDATA,
    output [32*6 -1: 0]     AXI_RID,
    output [32*1-1:0]   AXI_RLAST,
    output [32*2 -1: 0]     AXI_RRESP,
    output [32*1-1:0]   AXI_RVALID,
    output [32*1-1:0]   AXI_WREADY,
    output [32*6 -1: 0]     AXI_BID,
    output [32*2 -1: 0]     AXI_BRESP,
    output [32*1-1:0]   AXI_BVALID,

    input hbm_diff_clk_p,
  
    input hbm_diff_clk_n

    // input axi_hbm_clk
);
  
  wire clk;
  wire HBM_REF_CLK_0;
  wire HBM_REF_CLK_1;
  wire  [31 : 0] APB_0_PWDATA;
  wire  [21 : 0] APB_0_PADDR;
  wire  APB_0_PCLK;
  wire  APB_0_PENABLE;
  wire  APB_0_PRESET_N;
  wire  APB_0_PSEL;
  wire  APB_0_PWRITE;
  wire  [31 : 0] APB_1_PWDATA;
  wire  [21 : 0] APB_1_PADDR;
  wire  APB_1_PCLK;
  wire  APB_1_PENABLE;
  wire  APB_1_PRESET_N;
  wire  APB_1_PSEL;
  wire  APB_1_PWRITE;

  assign APB_0_PWDATA=0;
  assign APB_0_PADDR=0;
  assign APB_0_PCLK=HBM_REF_CLK_0;
  assign APB_0_PENABLE=0;
  assign APB_0_PRESET_N=1;
  assign APB_0_PSEL=0;
  assign APB_0_PWRITE=0;

  assign APB_1_PWDATA=0;
  assign APB_1_PADDR=0;
  assign APB_1_PCLK=HBM_REF_CLK_0;
  assign APB_1_PENABLE=0;
  assign APB_1_PRESET_N=1;
  assign APB_1_PSEL=0;
  assign APB_1_PWRITE=0;

  assign HBM_REF_CLK_0 = clk;
  assign HBM_REF_CLK_1 = clk;

    hbm_clk_wiz hbm_clk_wiz
   (
    // Clock out ports
    .clk_out1(clk),     // output clk_out1
   // Clock in ports
    .clk_in1_p(hbm_diff_clk_p),    // input clk_in1_p
    .clk_in1_n(hbm_diff_clk_n)    // input clk_in1_n
);

    hbm_0 hbm (
  .HBM_REF_CLK_0(HBM_REF_CLK_0),              // input wire HBM_REF_CLK_0
  .HBM_REF_CLK_1(HBM_REF_CLK_1),              // input wire HBM_REF_CLK_1

    .AXI_00_ACLK(AXI_ACLK[`getvec(1,0)]),
    .AXI_00_ARESET_N(AXI_ARESET_N[`getvec(1,0)]),
    .AXI_00_ARADDR(AXI_ARADDR[`getvec(33,0)]),
    .AXI_00_ARBURST(AXI_ARBURST[`getvec(2,0)]),
    .AXI_00_ARID(AXI_ARID[`getvec(6,0)]),
    .AXI_00_ARLEN(AXI_ARLEN[`getvec(4,0)]),
    .AXI_00_ARSIZE(AXI_ARSIZE[`getvec(3,0)]),
    .AXI_00_ARVALID(AXI_ARVALID[`getvec(1,0)]),
    .AXI_00_AWADDR(AXI_AWADDR[`getvec(33,0)]),
    .AXI_00_AWBURST(AXI_AWBURST[`getvec(2,0)]),
    .AXI_00_AWID(AXI_AWID[`getvec(6,0)]),
    .AXI_00_AWLEN(AXI_AWLEN[`getvec(4,0)]),
    .AXI_00_AWSIZE(AXI_AWSIZE[`getvec(3,0)]),
    .AXI_00_AWVALID(AXI_AWVALID[`getvec(1,0)]),
    .AXI_00_RREADY(AXI_RREADY[`getvec(1,0)]),
    .AXI_00_BREADY(AXI_BREADY[`getvec(1,0)]),
    .AXI_00_WDATA(AXI_WDATA[`getvec(256,0)]),
    .AXI_00_WLAST(AXI_WLAST[`getvec(1,0)]),
    .AXI_00_WSTRB(AXI_WSTRB[`getvec(32,0)]),
    .AXI_00_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,0)]),
    .AXI_00_WVALID(AXI_WVALID[`getvec(1,0)]),
    .AXI_00_ARREADY(AXI_ARREADY[`getvec(1,0)]),
    .AXI_00_AWREADY(AXI_AWREADY[`getvec(1,0)]),
    .AXI_00_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,0)]),
    .AXI_00_RDATA(AXI_RDATA[`getvec(256,0)]),
    .AXI_00_RID(AXI_RID[`getvec(6,0)]),
    .AXI_00_RLAST(AXI_RLAST[`getvec(1,0)]),
    .AXI_00_RRESP(AXI_RRESP[`getvec(2,0)]),
    .AXI_00_RVALID(AXI_RVALID[`getvec(1,0)]),
    .AXI_00_WREADY(AXI_WREADY[`getvec(1,0)]),
    .AXI_00_BID(AXI_BID[`getvec(6,0)]),
    .AXI_00_BRESP(AXI_BRESP[`getvec(2,0)]),
    .AXI_00_BVALID(AXI_BVALID[`getvec(1,0)]),
    .AXI_01_ACLK(AXI_ACLK[`getvec(1,1)]),
    .AXI_01_ARESET_N(AXI_ARESET_N[`getvec(1,1)]),
    .AXI_01_ARADDR(AXI_ARADDR[`getvec(33,1)]),
    .AXI_01_ARBURST(AXI_ARBURST[`getvec(2,1)]),
    .AXI_01_ARID(AXI_ARID[`getvec(6,1)]),
    .AXI_01_ARLEN(AXI_ARLEN[`getvec(4,1)]),
    .AXI_01_ARSIZE(AXI_ARSIZE[`getvec(3,1)]),
    .AXI_01_ARVALID(AXI_ARVALID[`getvec(1,1)]),
    .AXI_01_AWADDR(AXI_AWADDR[`getvec(33,1)]),
    .AXI_01_AWBURST(AXI_AWBURST[`getvec(2,1)]),
    .AXI_01_AWID(AXI_AWID[`getvec(6,1)]),
    .AXI_01_AWLEN(AXI_AWLEN[`getvec(4,1)]),
    .AXI_01_AWSIZE(AXI_AWSIZE[`getvec(3,1)]),
    .AXI_01_AWVALID(AXI_AWVALID[`getvec(1,1)]),
    .AXI_01_RREADY(AXI_RREADY[`getvec(1,1)]),
    .AXI_01_BREADY(AXI_BREADY[`getvec(1,1)]),
    .AXI_01_WDATA(AXI_WDATA[`getvec(256,1)]),
    .AXI_01_WLAST(AXI_WLAST[`getvec(1,1)]),
    .AXI_01_WSTRB(AXI_WSTRB[`getvec(32,1)]),
    .AXI_01_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,1)]),
    .AXI_01_WVALID(AXI_WVALID[`getvec(1,1)]),
    .AXI_01_ARREADY(AXI_ARREADY[`getvec(1,1)]),
    .AXI_01_AWREADY(AXI_AWREADY[`getvec(1,1)]),
    .AXI_01_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,1)]),
    .AXI_01_RDATA(AXI_RDATA[`getvec(256,1)]),
    .AXI_01_RID(AXI_RID[`getvec(6,1)]),
    .AXI_01_RLAST(AXI_RLAST[`getvec(1,1)]),
    .AXI_01_RRESP(AXI_RRESP[`getvec(2,1)]),
    .AXI_01_RVALID(AXI_RVALID[`getvec(1,1)]),
    .AXI_01_WREADY(AXI_WREADY[`getvec(1,1)]),
    .AXI_01_BID(AXI_BID[`getvec(6,1)]),
    .AXI_01_BRESP(AXI_BRESP[`getvec(2,1)]),
    .AXI_01_BVALID(AXI_BVALID[`getvec(1,1)]),
    .AXI_02_ACLK(AXI_ACLK[`getvec(1,2)]),
    .AXI_02_ARESET_N(AXI_ARESET_N[`getvec(1,2)]),
    .AXI_02_ARADDR(AXI_ARADDR[`getvec(33,2)]),
    .AXI_02_ARBURST(AXI_ARBURST[`getvec(2,2)]),
    .AXI_02_ARID(AXI_ARID[`getvec(6,2)]),
    .AXI_02_ARLEN(AXI_ARLEN[`getvec(4,2)]),
    .AXI_02_ARSIZE(AXI_ARSIZE[`getvec(3,2)]),
    .AXI_02_ARVALID(AXI_ARVALID[`getvec(1,2)]),
    .AXI_02_AWADDR(AXI_AWADDR[`getvec(33,2)]),
    .AXI_02_AWBURST(AXI_AWBURST[`getvec(2,2)]),
    .AXI_02_AWID(AXI_AWID[`getvec(6,2)]),
    .AXI_02_AWLEN(AXI_AWLEN[`getvec(4,2)]),
    .AXI_02_AWSIZE(AXI_AWSIZE[`getvec(3,2)]),
    .AXI_02_AWVALID(AXI_AWVALID[`getvec(1,2)]),
    .AXI_02_RREADY(AXI_RREADY[`getvec(1,2)]),
    .AXI_02_BREADY(AXI_BREADY[`getvec(1,2)]),
    .AXI_02_WDATA(AXI_WDATA[`getvec(256,2)]),
    .AXI_02_WLAST(AXI_WLAST[`getvec(1,2)]),
    .AXI_02_WSTRB(AXI_WSTRB[`getvec(32,2)]),
    .AXI_02_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,2)]),
    .AXI_02_WVALID(AXI_WVALID[`getvec(1,2)]),
    .AXI_02_ARREADY(AXI_ARREADY[`getvec(1,2)]),
    .AXI_02_AWREADY(AXI_AWREADY[`getvec(1,2)]),
    .AXI_02_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,2)]),
    .AXI_02_RDATA(AXI_RDATA[`getvec(256,2)]),
    .AXI_02_RID(AXI_RID[`getvec(6,2)]),
    .AXI_02_RLAST(AXI_RLAST[`getvec(1,2)]),
    .AXI_02_RRESP(AXI_RRESP[`getvec(2,2)]),
    .AXI_02_RVALID(AXI_RVALID[`getvec(1,2)]),
    .AXI_02_WREADY(AXI_WREADY[`getvec(1,2)]),
    .AXI_02_BID(AXI_BID[`getvec(6,2)]),
    .AXI_02_BRESP(AXI_BRESP[`getvec(2,2)]),
    .AXI_02_BVALID(AXI_BVALID[`getvec(1,2)]),
    .AXI_03_ACLK(AXI_ACLK[`getvec(1,3)]),
    .AXI_03_ARESET_N(AXI_ARESET_N[`getvec(1,3)]),
    .AXI_03_ARADDR(AXI_ARADDR[`getvec(33,3)]),
    .AXI_03_ARBURST(AXI_ARBURST[`getvec(2,3)]),
    .AXI_03_ARID(AXI_ARID[`getvec(6,3)]),
    .AXI_03_ARLEN(AXI_ARLEN[`getvec(4,3)]),
    .AXI_03_ARSIZE(AXI_ARSIZE[`getvec(3,3)]),
    .AXI_03_ARVALID(AXI_ARVALID[`getvec(1,3)]),
    .AXI_03_AWADDR(AXI_AWADDR[`getvec(33,3)]),
    .AXI_03_AWBURST(AXI_AWBURST[`getvec(2,3)]),
    .AXI_03_AWID(AXI_AWID[`getvec(6,3)]),
    .AXI_03_AWLEN(AXI_AWLEN[`getvec(4,3)]),
    .AXI_03_AWSIZE(AXI_AWSIZE[`getvec(3,3)]),
    .AXI_03_AWVALID(AXI_AWVALID[`getvec(1,3)]),
    .AXI_03_RREADY(AXI_RREADY[`getvec(1,3)]),
    .AXI_03_BREADY(AXI_BREADY[`getvec(1,3)]),
    .AXI_03_WDATA(AXI_WDATA[`getvec(256,3)]),
    .AXI_03_WLAST(AXI_WLAST[`getvec(1,3)]),
    .AXI_03_WSTRB(AXI_WSTRB[`getvec(32,3)]),
    .AXI_03_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,3)]),
    .AXI_03_WVALID(AXI_WVALID[`getvec(1,3)]),
    .AXI_03_ARREADY(AXI_ARREADY[`getvec(1,3)]),
    .AXI_03_AWREADY(AXI_AWREADY[`getvec(1,3)]),
    .AXI_03_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,3)]),
    .AXI_03_RDATA(AXI_RDATA[`getvec(256,3)]),
    .AXI_03_RID(AXI_RID[`getvec(6,3)]),
    .AXI_03_RLAST(AXI_RLAST[`getvec(1,3)]),
    .AXI_03_RRESP(AXI_RRESP[`getvec(2,3)]),
    .AXI_03_RVALID(AXI_RVALID[`getvec(1,3)]),
    .AXI_03_WREADY(AXI_WREADY[`getvec(1,3)]),
    .AXI_03_BID(AXI_BID[`getvec(6,3)]),
    .AXI_03_BRESP(AXI_BRESP[`getvec(2,3)]),
    .AXI_03_BVALID(AXI_BVALID[`getvec(1,3)]),
    .AXI_04_ACLK(AXI_ACLK[`getvec(1,4)]),
    .AXI_04_ARESET_N(AXI_ARESET_N[`getvec(1,4)]),
    .AXI_04_ARADDR(AXI_ARADDR[`getvec(33,4)]),
    .AXI_04_ARBURST(AXI_ARBURST[`getvec(2,4)]),
    .AXI_04_ARID(AXI_ARID[`getvec(6,4)]),
    .AXI_04_ARLEN(AXI_ARLEN[`getvec(4,4)]),
    .AXI_04_ARSIZE(AXI_ARSIZE[`getvec(3,4)]),
    .AXI_04_ARVALID(AXI_ARVALID[`getvec(1,4)]),
    .AXI_04_AWADDR(AXI_AWADDR[`getvec(33,4)]),
    .AXI_04_AWBURST(AXI_AWBURST[`getvec(2,4)]),
    .AXI_04_AWID(AXI_AWID[`getvec(6,4)]),
    .AXI_04_AWLEN(AXI_AWLEN[`getvec(4,4)]),
    .AXI_04_AWSIZE(AXI_AWSIZE[`getvec(3,4)]),
    .AXI_04_AWVALID(AXI_AWVALID[`getvec(1,4)]),
    .AXI_04_RREADY(AXI_RREADY[`getvec(1,4)]),
    .AXI_04_BREADY(AXI_BREADY[`getvec(1,4)]),
    .AXI_04_WDATA(AXI_WDATA[`getvec(256,4)]),
    .AXI_04_WLAST(AXI_WLAST[`getvec(1,4)]),
    .AXI_04_WSTRB(AXI_WSTRB[`getvec(32,4)]),
    .AXI_04_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,4)]),
    .AXI_04_WVALID(AXI_WVALID[`getvec(1,4)]),
    .AXI_04_ARREADY(AXI_ARREADY[`getvec(1,4)]),
    .AXI_04_AWREADY(AXI_AWREADY[`getvec(1,4)]),
    .AXI_04_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,4)]),
    .AXI_04_RDATA(AXI_RDATA[`getvec(256,4)]),
    .AXI_04_RID(AXI_RID[`getvec(6,4)]),
    .AXI_04_RLAST(AXI_RLAST[`getvec(1,4)]),
    .AXI_04_RRESP(AXI_RRESP[`getvec(2,4)]),
    .AXI_04_RVALID(AXI_RVALID[`getvec(1,4)]),
    .AXI_04_WREADY(AXI_WREADY[`getvec(1,4)]),
    .AXI_04_BID(AXI_BID[`getvec(6,4)]),
    .AXI_04_BRESP(AXI_BRESP[`getvec(2,4)]),
    .AXI_04_BVALID(AXI_BVALID[`getvec(1,4)]),
    .AXI_05_ACLK(AXI_ACLK[`getvec(1,5)]),
    .AXI_05_ARESET_N(AXI_ARESET_N[`getvec(1,5)]),
    .AXI_05_ARADDR(AXI_ARADDR[`getvec(33,5)]),
    .AXI_05_ARBURST(AXI_ARBURST[`getvec(2,5)]),
    .AXI_05_ARID(AXI_ARID[`getvec(6,5)]),
    .AXI_05_ARLEN(AXI_ARLEN[`getvec(4,5)]),
    .AXI_05_ARSIZE(AXI_ARSIZE[`getvec(3,5)]),
    .AXI_05_ARVALID(AXI_ARVALID[`getvec(1,5)]),
    .AXI_05_AWADDR(AXI_AWADDR[`getvec(33,5)]),
    .AXI_05_AWBURST(AXI_AWBURST[`getvec(2,5)]),
    .AXI_05_AWID(AXI_AWID[`getvec(6,5)]),
    .AXI_05_AWLEN(AXI_AWLEN[`getvec(4,5)]),
    .AXI_05_AWSIZE(AXI_AWSIZE[`getvec(3,5)]),
    .AXI_05_AWVALID(AXI_AWVALID[`getvec(1,5)]),
    .AXI_05_RREADY(AXI_RREADY[`getvec(1,5)]),
    .AXI_05_BREADY(AXI_BREADY[`getvec(1,5)]),
    .AXI_05_WDATA(AXI_WDATA[`getvec(256,5)]),
    .AXI_05_WLAST(AXI_WLAST[`getvec(1,5)]),
    .AXI_05_WSTRB(AXI_WSTRB[`getvec(32,5)]),
    .AXI_05_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,5)]),
    .AXI_05_WVALID(AXI_WVALID[`getvec(1,5)]),
    .AXI_05_ARREADY(AXI_ARREADY[`getvec(1,5)]),
    .AXI_05_AWREADY(AXI_AWREADY[`getvec(1,5)]),
    .AXI_05_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,5)]),
    .AXI_05_RDATA(AXI_RDATA[`getvec(256,5)]),
    .AXI_05_RID(AXI_RID[`getvec(6,5)]),
    .AXI_05_RLAST(AXI_RLAST[`getvec(1,5)]),
    .AXI_05_RRESP(AXI_RRESP[`getvec(2,5)]),
    .AXI_05_RVALID(AXI_RVALID[`getvec(1,5)]),
    .AXI_05_WREADY(AXI_WREADY[`getvec(1,5)]),
    .AXI_05_BID(AXI_BID[`getvec(6,5)]),
    .AXI_05_BRESP(AXI_BRESP[`getvec(2,5)]),
    .AXI_05_BVALID(AXI_BVALID[`getvec(1,5)]),
    .AXI_06_ACLK(AXI_ACLK[`getvec(1,6)]),
    .AXI_06_ARESET_N(AXI_ARESET_N[`getvec(1,6)]),
    .AXI_06_ARADDR(AXI_ARADDR[`getvec(33,6)]),
    .AXI_06_ARBURST(AXI_ARBURST[`getvec(2,6)]),
    .AXI_06_ARID(AXI_ARID[`getvec(6,6)]),
    .AXI_06_ARLEN(AXI_ARLEN[`getvec(4,6)]),
    .AXI_06_ARSIZE(AXI_ARSIZE[`getvec(3,6)]),
    .AXI_06_ARVALID(AXI_ARVALID[`getvec(1,6)]),
    .AXI_06_AWADDR(AXI_AWADDR[`getvec(33,6)]),
    .AXI_06_AWBURST(AXI_AWBURST[`getvec(2,6)]),
    .AXI_06_AWID(AXI_AWID[`getvec(6,6)]),
    .AXI_06_AWLEN(AXI_AWLEN[`getvec(4,6)]),
    .AXI_06_AWSIZE(AXI_AWSIZE[`getvec(3,6)]),
    .AXI_06_AWVALID(AXI_AWVALID[`getvec(1,6)]),
    .AXI_06_RREADY(AXI_RREADY[`getvec(1,6)]),
    .AXI_06_BREADY(AXI_BREADY[`getvec(1,6)]),
    .AXI_06_WDATA(AXI_WDATA[`getvec(256,6)]),
    .AXI_06_WLAST(AXI_WLAST[`getvec(1,6)]),
    .AXI_06_WSTRB(AXI_WSTRB[`getvec(32,6)]),
    .AXI_06_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,6)]),
    .AXI_06_WVALID(AXI_WVALID[`getvec(1,6)]),
    .AXI_06_ARREADY(AXI_ARREADY[`getvec(1,6)]),
    .AXI_06_AWREADY(AXI_AWREADY[`getvec(1,6)]),
    .AXI_06_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,6)]),
    .AXI_06_RDATA(AXI_RDATA[`getvec(256,6)]),
    .AXI_06_RID(AXI_RID[`getvec(6,6)]),
    .AXI_06_RLAST(AXI_RLAST[`getvec(1,6)]),
    .AXI_06_RRESP(AXI_RRESP[`getvec(2,6)]),
    .AXI_06_RVALID(AXI_RVALID[`getvec(1,6)]),
    .AXI_06_WREADY(AXI_WREADY[`getvec(1,6)]),
    .AXI_06_BID(AXI_BID[`getvec(6,6)]),
    .AXI_06_BRESP(AXI_BRESP[`getvec(2,6)]),
    .AXI_06_BVALID(AXI_BVALID[`getvec(1,6)]),
    .AXI_07_ACLK(AXI_ACLK[`getvec(1,7)]),
    .AXI_07_ARESET_N(AXI_ARESET_N[`getvec(1,7)]),
    .AXI_07_ARADDR(AXI_ARADDR[`getvec(33,7)]),
    .AXI_07_ARBURST(AXI_ARBURST[`getvec(2,7)]),
    .AXI_07_ARID(AXI_ARID[`getvec(6,7)]),
    .AXI_07_ARLEN(AXI_ARLEN[`getvec(4,7)]),
    .AXI_07_ARSIZE(AXI_ARSIZE[`getvec(3,7)]),
    .AXI_07_ARVALID(AXI_ARVALID[`getvec(1,7)]),
    .AXI_07_AWADDR(AXI_AWADDR[`getvec(33,7)]),
    .AXI_07_AWBURST(AXI_AWBURST[`getvec(2,7)]),
    .AXI_07_AWID(AXI_AWID[`getvec(6,7)]),
    .AXI_07_AWLEN(AXI_AWLEN[`getvec(4,7)]),
    .AXI_07_AWSIZE(AXI_AWSIZE[`getvec(3,7)]),
    .AXI_07_AWVALID(AXI_AWVALID[`getvec(1,7)]),
    .AXI_07_RREADY(AXI_RREADY[`getvec(1,7)]),
    .AXI_07_BREADY(AXI_BREADY[`getvec(1,7)]),
    .AXI_07_WDATA(AXI_WDATA[`getvec(256,7)]),
    .AXI_07_WLAST(AXI_WLAST[`getvec(1,7)]),
    .AXI_07_WSTRB(AXI_WSTRB[`getvec(32,7)]),
    .AXI_07_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,7)]),
    .AXI_07_WVALID(AXI_WVALID[`getvec(1,7)]),
    .AXI_07_ARREADY(AXI_ARREADY[`getvec(1,7)]),
    .AXI_07_AWREADY(AXI_AWREADY[`getvec(1,7)]),
    .AXI_07_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,7)]),
    .AXI_07_RDATA(AXI_RDATA[`getvec(256,7)]),
    .AXI_07_RID(AXI_RID[`getvec(6,7)]),
    .AXI_07_RLAST(AXI_RLAST[`getvec(1,7)]),
    .AXI_07_RRESP(AXI_RRESP[`getvec(2,7)]),
    .AXI_07_RVALID(AXI_RVALID[`getvec(1,7)]),
    .AXI_07_WREADY(AXI_WREADY[`getvec(1,7)]),
    .AXI_07_BID(AXI_BID[`getvec(6,7)]),
    .AXI_07_BRESP(AXI_BRESP[`getvec(2,7)]),
    .AXI_07_BVALID(AXI_BVALID[`getvec(1,7)]),
    .AXI_08_ACLK(AXI_ACLK[`getvec(1,8)]),
    .AXI_08_ARESET_N(AXI_ARESET_N[`getvec(1,8)]),
    .AXI_08_ARADDR(AXI_ARADDR[`getvec(33,8)]),
    .AXI_08_ARBURST(AXI_ARBURST[`getvec(2,8)]),
    .AXI_08_ARID(AXI_ARID[`getvec(6,8)]),
    .AXI_08_ARLEN(AXI_ARLEN[`getvec(4,8)]),
    .AXI_08_ARSIZE(AXI_ARSIZE[`getvec(3,8)]),
    .AXI_08_ARVALID(AXI_ARVALID[`getvec(1,8)]),
    .AXI_08_AWADDR(AXI_AWADDR[`getvec(33,8)]),
    .AXI_08_AWBURST(AXI_AWBURST[`getvec(2,8)]),
    .AXI_08_AWID(AXI_AWID[`getvec(6,8)]),
    .AXI_08_AWLEN(AXI_AWLEN[`getvec(4,8)]),
    .AXI_08_AWSIZE(AXI_AWSIZE[`getvec(3,8)]),
    .AXI_08_AWVALID(AXI_AWVALID[`getvec(1,8)]),
    .AXI_08_RREADY(AXI_RREADY[`getvec(1,8)]),
    .AXI_08_BREADY(AXI_BREADY[`getvec(1,8)]),
    .AXI_08_WDATA(AXI_WDATA[`getvec(256,8)]),
    .AXI_08_WLAST(AXI_WLAST[`getvec(1,8)]),
    .AXI_08_WSTRB(AXI_WSTRB[`getvec(32,8)]),
    .AXI_08_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,8)]),
    .AXI_08_WVALID(AXI_WVALID[`getvec(1,8)]),
    .AXI_08_ARREADY(AXI_ARREADY[`getvec(1,8)]),
    .AXI_08_AWREADY(AXI_AWREADY[`getvec(1,8)]),
    .AXI_08_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,8)]),
    .AXI_08_RDATA(AXI_RDATA[`getvec(256,8)]),
    .AXI_08_RID(AXI_RID[`getvec(6,8)]),
    .AXI_08_RLAST(AXI_RLAST[`getvec(1,8)]),
    .AXI_08_RRESP(AXI_RRESP[`getvec(2,8)]),
    .AXI_08_RVALID(AXI_RVALID[`getvec(1,8)]),
    .AXI_08_WREADY(AXI_WREADY[`getvec(1,8)]),
    .AXI_08_BID(AXI_BID[`getvec(6,8)]),
    .AXI_08_BRESP(AXI_BRESP[`getvec(2,8)]),
    .AXI_08_BVALID(AXI_BVALID[`getvec(1,8)]),
    .AXI_09_ACLK(AXI_ACLK[`getvec(1,9)]),
    .AXI_09_ARESET_N(AXI_ARESET_N[`getvec(1,9)]),
    .AXI_09_ARADDR(AXI_ARADDR[`getvec(33,9)]),
    .AXI_09_ARBURST(AXI_ARBURST[`getvec(2,9)]),
    .AXI_09_ARID(AXI_ARID[`getvec(6,9)]),
    .AXI_09_ARLEN(AXI_ARLEN[`getvec(4,9)]),
    .AXI_09_ARSIZE(AXI_ARSIZE[`getvec(3,9)]),
    .AXI_09_ARVALID(AXI_ARVALID[`getvec(1,9)]),
    .AXI_09_AWADDR(AXI_AWADDR[`getvec(33,9)]),
    .AXI_09_AWBURST(AXI_AWBURST[`getvec(2,9)]),
    .AXI_09_AWID(AXI_AWID[`getvec(6,9)]),
    .AXI_09_AWLEN(AXI_AWLEN[`getvec(4,9)]),
    .AXI_09_AWSIZE(AXI_AWSIZE[`getvec(3,9)]),
    .AXI_09_AWVALID(AXI_AWVALID[`getvec(1,9)]),
    .AXI_09_RREADY(AXI_RREADY[`getvec(1,9)]),
    .AXI_09_BREADY(AXI_BREADY[`getvec(1,9)]),
    .AXI_09_WDATA(AXI_WDATA[`getvec(256,9)]),
    .AXI_09_WLAST(AXI_WLAST[`getvec(1,9)]),
    .AXI_09_WSTRB(AXI_WSTRB[`getvec(32,9)]),
    .AXI_09_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,9)]),
    .AXI_09_WVALID(AXI_WVALID[`getvec(1,9)]),
    .AXI_09_ARREADY(AXI_ARREADY[`getvec(1,9)]),
    .AXI_09_AWREADY(AXI_AWREADY[`getvec(1,9)]),
    .AXI_09_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,9)]),
    .AXI_09_RDATA(AXI_RDATA[`getvec(256,9)]),
    .AXI_09_RID(AXI_RID[`getvec(6,9)]),
    .AXI_09_RLAST(AXI_RLAST[`getvec(1,9)]),
    .AXI_09_RRESP(AXI_RRESP[`getvec(2,9)]),
    .AXI_09_RVALID(AXI_RVALID[`getvec(1,9)]),
    .AXI_09_WREADY(AXI_WREADY[`getvec(1,9)]),
    .AXI_09_BID(AXI_BID[`getvec(6,9)]),
    .AXI_09_BRESP(AXI_BRESP[`getvec(2,9)]),
    .AXI_09_BVALID(AXI_BVALID[`getvec(1,9)]),
    .AXI_10_ACLK(AXI_ACLK[`getvec(1,10)]),
    .AXI_10_ARESET_N(AXI_ARESET_N[`getvec(1,10)]),
    .AXI_10_ARADDR(AXI_ARADDR[`getvec(33,10)]),
    .AXI_10_ARBURST(AXI_ARBURST[`getvec(2,10)]),
    .AXI_10_ARID(AXI_ARID[`getvec(6,10)]),
    .AXI_10_ARLEN(AXI_ARLEN[`getvec(4,10)]),
    .AXI_10_ARSIZE(AXI_ARSIZE[`getvec(3,10)]),
    .AXI_10_ARVALID(AXI_ARVALID[`getvec(1,10)]),
    .AXI_10_AWADDR(AXI_AWADDR[`getvec(33,10)]),
    .AXI_10_AWBURST(AXI_AWBURST[`getvec(2,10)]),
    .AXI_10_AWID(AXI_AWID[`getvec(6,10)]),
    .AXI_10_AWLEN(AXI_AWLEN[`getvec(4,10)]),
    .AXI_10_AWSIZE(AXI_AWSIZE[`getvec(3,10)]),
    .AXI_10_AWVALID(AXI_AWVALID[`getvec(1,10)]),
    .AXI_10_RREADY(AXI_RREADY[`getvec(1,10)]),
    .AXI_10_BREADY(AXI_BREADY[`getvec(1,10)]),
    .AXI_10_WDATA(AXI_WDATA[`getvec(256,10)]),
    .AXI_10_WLAST(AXI_WLAST[`getvec(1,10)]),
    .AXI_10_WSTRB(AXI_WSTRB[`getvec(32,10)]),
    .AXI_10_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,10)]),
    .AXI_10_WVALID(AXI_WVALID[`getvec(1,10)]),
    .AXI_10_ARREADY(AXI_ARREADY[`getvec(1,10)]),
    .AXI_10_AWREADY(AXI_AWREADY[`getvec(1,10)]),
    .AXI_10_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,10)]),
    .AXI_10_RDATA(AXI_RDATA[`getvec(256,10)]),
    .AXI_10_RID(AXI_RID[`getvec(6,10)]),
    .AXI_10_RLAST(AXI_RLAST[`getvec(1,10)]),
    .AXI_10_RRESP(AXI_RRESP[`getvec(2,10)]),
    .AXI_10_RVALID(AXI_RVALID[`getvec(1,10)]),
    .AXI_10_WREADY(AXI_WREADY[`getvec(1,10)]),
    .AXI_10_BID(AXI_BID[`getvec(6,10)]),
    .AXI_10_BRESP(AXI_BRESP[`getvec(2,10)]),
    .AXI_10_BVALID(AXI_BVALID[`getvec(1,10)]),
    .AXI_11_ACLK(AXI_ACLK[`getvec(1,11)]),
    .AXI_11_ARESET_N(AXI_ARESET_N[`getvec(1,11)]),
    .AXI_11_ARADDR(AXI_ARADDR[`getvec(33,11)]),
    .AXI_11_ARBURST(AXI_ARBURST[`getvec(2,11)]),
    .AXI_11_ARID(AXI_ARID[`getvec(6,11)]),
    .AXI_11_ARLEN(AXI_ARLEN[`getvec(4,11)]),
    .AXI_11_ARSIZE(AXI_ARSIZE[`getvec(3,11)]),
    .AXI_11_ARVALID(AXI_ARVALID[`getvec(1,11)]),
    .AXI_11_AWADDR(AXI_AWADDR[`getvec(33,11)]),
    .AXI_11_AWBURST(AXI_AWBURST[`getvec(2,11)]),
    .AXI_11_AWID(AXI_AWID[`getvec(6,11)]),
    .AXI_11_AWLEN(AXI_AWLEN[`getvec(4,11)]),
    .AXI_11_AWSIZE(AXI_AWSIZE[`getvec(3,11)]),
    .AXI_11_AWVALID(AXI_AWVALID[`getvec(1,11)]),
    .AXI_11_RREADY(AXI_RREADY[`getvec(1,11)]),
    .AXI_11_BREADY(AXI_BREADY[`getvec(1,11)]),
    .AXI_11_WDATA(AXI_WDATA[`getvec(256,11)]),
    .AXI_11_WLAST(AXI_WLAST[`getvec(1,11)]),
    .AXI_11_WSTRB(AXI_WSTRB[`getvec(32,11)]),
    .AXI_11_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,11)]),
    .AXI_11_WVALID(AXI_WVALID[`getvec(1,11)]),
    .AXI_11_ARREADY(AXI_ARREADY[`getvec(1,11)]),
    .AXI_11_AWREADY(AXI_AWREADY[`getvec(1,11)]),
    .AXI_11_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,11)]),
    .AXI_11_RDATA(AXI_RDATA[`getvec(256,11)]),
    .AXI_11_RID(AXI_RID[`getvec(6,11)]),
    .AXI_11_RLAST(AXI_RLAST[`getvec(1,11)]),
    .AXI_11_RRESP(AXI_RRESP[`getvec(2,11)]),
    .AXI_11_RVALID(AXI_RVALID[`getvec(1,11)]),
    .AXI_11_WREADY(AXI_WREADY[`getvec(1,11)]),
    .AXI_11_BID(AXI_BID[`getvec(6,11)]),
    .AXI_11_BRESP(AXI_BRESP[`getvec(2,11)]),
    .AXI_11_BVALID(AXI_BVALID[`getvec(1,11)]),
    .AXI_12_ACLK(AXI_ACLK[`getvec(1,12)]),
    .AXI_12_ARESET_N(AXI_ARESET_N[`getvec(1,12)]),
    .AXI_12_ARADDR(AXI_ARADDR[`getvec(33,12)]),
    .AXI_12_ARBURST(AXI_ARBURST[`getvec(2,12)]),
    .AXI_12_ARID(AXI_ARID[`getvec(6,12)]),
    .AXI_12_ARLEN(AXI_ARLEN[`getvec(4,12)]),
    .AXI_12_ARSIZE(AXI_ARSIZE[`getvec(3,12)]),
    .AXI_12_ARVALID(AXI_ARVALID[`getvec(1,12)]),
    .AXI_12_AWADDR(AXI_AWADDR[`getvec(33,12)]),
    .AXI_12_AWBURST(AXI_AWBURST[`getvec(2,12)]),
    .AXI_12_AWID(AXI_AWID[`getvec(6,12)]),
    .AXI_12_AWLEN(AXI_AWLEN[`getvec(4,12)]),
    .AXI_12_AWSIZE(AXI_AWSIZE[`getvec(3,12)]),
    .AXI_12_AWVALID(AXI_AWVALID[`getvec(1,12)]),
    .AXI_12_RREADY(AXI_RREADY[`getvec(1,12)]),
    .AXI_12_BREADY(AXI_BREADY[`getvec(1,12)]),
    .AXI_12_WDATA(AXI_WDATA[`getvec(256,12)]),
    .AXI_12_WLAST(AXI_WLAST[`getvec(1,12)]),
    .AXI_12_WSTRB(AXI_WSTRB[`getvec(32,12)]),
    .AXI_12_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,12)]),
    .AXI_12_WVALID(AXI_WVALID[`getvec(1,12)]),
    .AXI_12_ARREADY(AXI_ARREADY[`getvec(1,12)]),
    .AXI_12_AWREADY(AXI_AWREADY[`getvec(1,12)]),
    .AXI_12_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,12)]),
    .AXI_12_RDATA(AXI_RDATA[`getvec(256,12)]),
    .AXI_12_RID(AXI_RID[`getvec(6,12)]),
    .AXI_12_RLAST(AXI_RLAST[`getvec(1,12)]),
    .AXI_12_RRESP(AXI_RRESP[`getvec(2,12)]),
    .AXI_12_RVALID(AXI_RVALID[`getvec(1,12)]),
    .AXI_12_WREADY(AXI_WREADY[`getvec(1,12)]),
    .AXI_12_BID(AXI_BID[`getvec(6,12)]),
    .AXI_12_BRESP(AXI_BRESP[`getvec(2,12)]),
    .AXI_12_BVALID(AXI_BVALID[`getvec(1,12)]),
    .AXI_13_ACLK(AXI_ACLK[`getvec(1,13)]),
    .AXI_13_ARESET_N(AXI_ARESET_N[`getvec(1,13)]),
    .AXI_13_ARADDR(AXI_ARADDR[`getvec(33,13)]),
    .AXI_13_ARBURST(AXI_ARBURST[`getvec(2,13)]),
    .AXI_13_ARID(AXI_ARID[`getvec(6,13)]),
    .AXI_13_ARLEN(AXI_ARLEN[`getvec(4,13)]),
    .AXI_13_ARSIZE(AXI_ARSIZE[`getvec(3,13)]),
    .AXI_13_ARVALID(AXI_ARVALID[`getvec(1,13)]),
    .AXI_13_AWADDR(AXI_AWADDR[`getvec(33,13)]),
    .AXI_13_AWBURST(AXI_AWBURST[`getvec(2,13)]),
    .AXI_13_AWID(AXI_AWID[`getvec(6,13)]),
    .AXI_13_AWLEN(AXI_AWLEN[`getvec(4,13)]),
    .AXI_13_AWSIZE(AXI_AWSIZE[`getvec(3,13)]),
    .AXI_13_AWVALID(AXI_AWVALID[`getvec(1,13)]),
    .AXI_13_RREADY(AXI_RREADY[`getvec(1,13)]),
    .AXI_13_BREADY(AXI_BREADY[`getvec(1,13)]),
    .AXI_13_WDATA(AXI_WDATA[`getvec(256,13)]),
    .AXI_13_WLAST(AXI_WLAST[`getvec(1,13)]),
    .AXI_13_WSTRB(AXI_WSTRB[`getvec(32,13)]),
    .AXI_13_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,13)]),
    .AXI_13_WVALID(AXI_WVALID[`getvec(1,13)]),
    .AXI_13_ARREADY(AXI_ARREADY[`getvec(1,13)]),
    .AXI_13_AWREADY(AXI_AWREADY[`getvec(1,13)]),
    .AXI_13_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,13)]),
    .AXI_13_RDATA(AXI_RDATA[`getvec(256,13)]),
    .AXI_13_RID(AXI_RID[`getvec(6,13)]),
    .AXI_13_RLAST(AXI_RLAST[`getvec(1,13)]),
    .AXI_13_RRESP(AXI_RRESP[`getvec(2,13)]),
    .AXI_13_RVALID(AXI_RVALID[`getvec(1,13)]),
    .AXI_13_WREADY(AXI_WREADY[`getvec(1,13)]),
    .AXI_13_BID(AXI_BID[`getvec(6,13)]),
    .AXI_13_BRESP(AXI_BRESP[`getvec(2,13)]),
    .AXI_13_BVALID(AXI_BVALID[`getvec(1,13)]),
    .AXI_14_ACLK(AXI_ACLK[`getvec(1,14)]),
    .AXI_14_ARESET_N(AXI_ARESET_N[`getvec(1,14)]),
    .AXI_14_ARADDR(AXI_ARADDR[`getvec(33,14)]),
    .AXI_14_ARBURST(AXI_ARBURST[`getvec(2,14)]),
    .AXI_14_ARID(AXI_ARID[`getvec(6,14)]),
    .AXI_14_ARLEN(AXI_ARLEN[`getvec(4,14)]),
    .AXI_14_ARSIZE(AXI_ARSIZE[`getvec(3,14)]),
    .AXI_14_ARVALID(AXI_ARVALID[`getvec(1,14)]),
    .AXI_14_AWADDR(AXI_AWADDR[`getvec(33,14)]),
    .AXI_14_AWBURST(AXI_AWBURST[`getvec(2,14)]),
    .AXI_14_AWID(AXI_AWID[`getvec(6,14)]),
    .AXI_14_AWLEN(AXI_AWLEN[`getvec(4,14)]),
    .AXI_14_AWSIZE(AXI_AWSIZE[`getvec(3,14)]),
    .AXI_14_AWVALID(AXI_AWVALID[`getvec(1,14)]),
    .AXI_14_RREADY(AXI_RREADY[`getvec(1,14)]),
    .AXI_14_BREADY(AXI_BREADY[`getvec(1,14)]),
    .AXI_14_WDATA(AXI_WDATA[`getvec(256,14)]),
    .AXI_14_WLAST(AXI_WLAST[`getvec(1,14)]),
    .AXI_14_WSTRB(AXI_WSTRB[`getvec(32,14)]),
    .AXI_14_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,14)]),
    .AXI_14_WVALID(AXI_WVALID[`getvec(1,14)]),
    .AXI_14_ARREADY(AXI_ARREADY[`getvec(1,14)]),
    .AXI_14_AWREADY(AXI_AWREADY[`getvec(1,14)]),
    .AXI_14_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,14)]),
    .AXI_14_RDATA(AXI_RDATA[`getvec(256,14)]),
    .AXI_14_RID(AXI_RID[`getvec(6,14)]),
    .AXI_14_RLAST(AXI_RLAST[`getvec(1,14)]),
    .AXI_14_RRESP(AXI_RRESP[`getvec(2,14)]),
    .AXI_14_RVALID(AXI_RVALID[`getvec(1,14)]),
    .AXI_14_WREADY(AXI_WREADY[`getvec(1,14)]),
    .AXI_14_BID(AXI_BID[`getvec(6,14)]),
    .AXI_14_BRESP(AXI_BRESP[`getvec(2,14)]),
    .AXI_14_BVALID(AXI_BVALID[`getvec(1,14)]),
    .AXI_15_ACLK(AXI_ACLK[`getvec(1,15)]),
    .AXI_15_ARESET_N(AXI_ARESET_N[`getvec(1,15)]),
    .AXI_15_ARADDR(AXI_ARADDR[`getvec(33,15)]),
    .AXI_15_ARBURST(AXI_ARBURST[`getvec(2,15)]),
    .AXI_15_ARID(AXI_ARID[`getvec(6,15)]),
    .AXI_15_ARLEN(AXI_ARLEN[`getvec(4,15)]),
    .AXI_15_ARSIZE(AXI_ARSIZE[`getvec(3,15)]),
    .AXI_15_ARVALID(AXI_ARVALID[`getvec(1,15)]),
    .AXI_15_AWADDR(AXI_AWADDR[`getvec(33,15)]),
    .AXI_15_AWBURST(AXI_AWBURST[`getvec(2,15)]),
    .AXI_15_AWID(AXI_AWID[`getvec(6,15)]),
    .AXI_15_AWLEN(AXI_AWLEN[`getvec(4,15)]),
    .AXI_15_AWSIZE(AXI_AWSIZE[`getvec(3,15)]),
    .AXI_15_AWVALID(AXI_AWVALID[`getvec(1,15)]),
    .AXI_15_RREADY(AXI_RREADY[`getvec(1,15)]),
    .AXI_15_BREADY(AXI_BREADY[`getvec(1,15)]),
    .AXI_15_WDATA(AXI_WDATA[`getvec(256,15)]),
    .AXI_15_WLAST(AXI_WLAST[`getvec(1,15)]),
    .AXI_15_WSTRB(AXI_WSTRB[`getvec(32,15)]),
    .AXI_15_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,15)]),
    .AXI_15_WVALID(AXI_WVALID[`getvec(1,15)]),
    .AXI_15_ARREADY(AXI_ARREADY[`getvec(1,15)]),
    .AXI_15_AWREADY(AXI_AWREADY[`getvec(1,15)]),
    .AXI_15_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,15)]),
    .AXI_15_RDATA(AXI_RDATA[`getvec(256,15)]),
    .AXI_15_RID(AXI_RID[`getvec(6,15)]),
    .AXI_15_RLAST(AXI_RLAST[`getvec(1,15)]),
    .AXI_15_RRESP(AXI_RRESP[`getvec(2,15)]),
    .AXI_15_RVALID(AXI_RVALID[`getvec(1,15)]),
    .AXI_15_WREADY(AXI_WREADY[`getvec(1,15)]),
    .AXI_15_BID(AXI_BID[`getvec(6,15)]),
    .AXI_15_BRESP(AXI_BRESP[`getvec(2,15)]),
    .AXI_15_BVALID(AXI_BVALID[`getvec(1,15)]),
    .AXI_16_ACLK(AXI_ACLK[`getvec(1,16)]),
    .AXI_16_ARESET_N(AXI_ARESET_N[`getvec(1,16)]),
    .AXI_16_ARADDR(AXI_ARADDR[`getvec(33,16)]),
    .AXI_16_ARBURST(AXI_ARBURST[`getvec(2,16)]),
    .AXI_16_ARID(AXI_ARID[`getvec(6,16)]),
    .AXI_16_ARLEN(AXI_ARLEN[`getvec(4,16)]),
    .AXI_16_ARSIZE(AXI_ARSIZE[`getvec(3,16)]),
    .AXI_16_ARVALID(AXI_ARVALID[`getvec(1,16)]),
    .AXI_16_AWADDR(AXI_AWADDR[`getvec(33,16)]),
    .AXI_16_AWBURST(AXI_AWBURST[`getvec(2,16)]),
    .AXI_16_AWID(AXI_AWID[`getvec(6,16)]),
    .AXI_16_AWLEN(AXI_AWLEN[`getvec(4,16)]),
    .AXI_16_AWSIZE(AXI_AWSIZE[`getvec(3,16)]),
    .AXI_16_AWVALID(AXI_AWVALID[`getvec(1,16)]),
    .AXI_16_RREADY(AXI_RREADY[`getvec(1,16)]),
    .AXI_16_BREADY(AXI_BREADY[`getvec(1,16)]),
    .AXI_16_WDATA(AXI_WDATA[`getvec(256,16)]),
    .AXI_16_WLAST(AXI_WLAST[`getvec(1,16)]),
    .AXI_16_WSTRB(AXI_WSTRB[`getvec(32,16)]),
    .AXI_16_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,16)]),
    .AXI_16_WVALID(AXI_WVALID[`getvec(1,16)]),
    .AXI_16_ARREADY(AXI_ARREADY[`getvec(1,16)]),
    .AXI_16_AWREADY(AXI_AWREADY[`getvec(1,16)]),
    .AXI_16_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,16)]),
    .AXI_16_RDATA(AXI_RDATA[`getvec(256,16)]),
    .AXI_16_RID(AXI_RID[`getvec(6,16)]),
    .AXI_16_RLAST(AXI_RLAST[`getvec(1,16)]),
    .AXI_16_RRESP(AXI_RRESP[`getvec(2,16)]),
    .AXI_16_RVALID(AXI_RVALID[`getvec(1,16)]),
    .AXI_16_WREADY(AXI_WREADY[`getvec(1,16)]),
    .AXI_16_BID(AXI_BID[`getvec(6,16)]),
    .AXI_16_BRESP(AXI_BRESP[`getvec(2,16)]),
    .AXI_16_BVALID(AXI_BVALID[`getvec(1,16)]),
    .AXI_17_ACLK(AXI_ACLK[`getvec(1,17)]),
    .AXI_17_ARESET_N(AXI_ARESET_N[`getvec(1,17)]),
    .AXI_17_ARADDR(AXI_ARADDR[`getvec(33,17)]),
    .AXI_17_ARBURST(AXI_ARBURST[`getvec(2,17)]),
    .AXI_17_ARID(AXI_ARID[`getvec(6,17)]),
    .AXI_17_ARLEN(AXI_ARLEN[`getvec(4,17)]),
    .AXI_17_ARSIZE(AXI_ARSIZE[`getvec(3,17)]),
    .AXI_17_ARVALID(AXI_ARVALID[`getvec(1,17)]),
    .AXI_17_AWADDR(AXI_AWADDR[`getvec(33,17)]),
    .AXI_17_AWBURST(AXI_AWBURST[`getvec(2,17)]),
    .AXI_17_AWID(AXI_AWID[`getvec(6,17)]),
    .AXI_17_AWLEN(AXI_AWLEN[`getvec(4,17)]),
    .AXI_17_AWSIZE(AXI_AWSIZE[`getvec(3,17)]),
    .AXI_17_AWVALID(AXI_AWVALID[`getvec(1,17)]),
    .AXI_17_RREADY(AXI_RREADY[`getvec(1,17)]),
    .AXI_17_BREADY(AXI_BREADY[`getvec(1,17)]),
    .AXI_17_WDATA(AXI_WDATA[`getvec(256,17)]),
    .AXI_17_WLAST(AXI_WLAST[`getvec(1,17)]),
    .AXI_17_WSTRB(AXI_WSTRB[`getvec(32,17)]),
    .AXI_17_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,17)]),
    .AXI_17_WVALID(AXI_WVALID[`getvec(1,17)]),
    .AXI_17_ARREADY(AXI_ARREADY[`getvec(1,17)]),
    .AXI_17_AWREADY(AXI_AWREADY[`getvec(1,17)]),
    .AXI_17_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,17)]),
    .AXI_17_RDATA(AXI_RDATA[`getvec(256,17)]),
    .AXI_17_RID(AXI_RID[`getvec(6,17)]),
    .AXI_17_RLAST(AXI_RLAST[`getvec(1,17)]),
    .AXI_17_RRESP(AXI_RRESP[`getvec(2,17)]),
    .AXI_17_RVALID(AXI_RVALID[`getvec(1,17)]),
    .AXI_17_WREADY(AXI_WREADY[`getvec(1,17)]),
    .AXI_17_BID(AXI_BID[`getvec(6,17)]),
    .AXI_17_BRESP(AXI_BRESP[`getvec(2,17)]),
    .AXI_17_BVALID(AXI_BVALID[`getvec(1,17)]),
    .AXI_18_ACLK(AXI_ACLK[`getvec(1,18)]),
    .AXI_18_ARESET_N(AXI_ARESET_N[`getvec(1,18)]),
    .AXI_18_ARADDR(AXI_ARADDR[`getvec(33,18)]),
    .AXI_18_ARBURST(AXI_ARBURST[`getvec(2,18)]),
    .AXI_18_ARID(AXI_ARID[`getvec(6,18)]),
    .AXI_18_ARLEN(AXI_ARLEN[`getvec(4,18)]),
    .AXI_18_ARSIZE(AXI_ARSIZE[`getvec(3,18)]),
    .AXI_18_ARVALID(AXI_ARVALID[`getvec(1,18)]),
    .AXI_18_AWADDR(AXI_AWADDR[`getvec(33,18)]),
    .AXI_18_AWBURST(AXI_AWBURST[`getvec(2,18)]),
    .AXI_18_AWID(AXI_AWID[`getvec(6,18)]),
    .AXI_18_AWLEN(AXI_AWLEN[`getvec(4,18)]),
    .AXI_18_AWSIZE(AXI_AWSIZE[`getvec(3,18)]),
    .AXI_18_AWVALID(AXI_AWVALID[`getvec(1,18)]),
    .AXI_18_RREADY(AXI_RREADY[`getvec(1,18)]),
    .AXI_18_BREADY(AXI_BREADY[`getvec(1,18)]),
    .AXI_18_WDATA(AXI_WDATA[`getvec(256,18)]),
    .AXI_18_WLAST(AXI_WLAST[`getvec(1,18)]),
    .AXI_18_WSTRB(AXI_WSTRB[`getvec(32,18)]),
    .AXI_18_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,18)]),
    .AXI_18_WVALID(AXI_WVALID[`getvec(1,18)]),
    .AXI_18_ARREADY(AXI_ARREADY[`getvec(1,18)]),
    .AXI_18_AWREADY(AXI_AWREADY[`getvec(1,18)]),
    .AXI_18_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,18)]),
    .AXI_18_RDATA(AXI_RDATA[`getvec(256,18)]),
    .AXI_18_RID(AXI_RID[`getvec(6,18)]),
    .AXI_18_RLAST(AXI_RLAST[`getvec(1,18)]),
    .AXI_18_RRESP(AXI_RRESP[`getvec(2,18)]),
    .AXI_18_RVALID(AXI_RVALID[`getvec(1,18)]),
    .AXI_18_WREADY(AXI_WREADY[`getvec(1,18)]),
    .AXI_18_BID(AXI_BID[`getvec(6,18)]),
    .AXI_18_BRESP(AXI_BRESP[`getvec(2,18)]),
    .AXI_18_BVALID(AXI_BVALID[`getvec(1,18)]),
    .AXI_19_ACLK(AXI_ACLK[`getvec(1,19)]),
    .AXI_19_ARESET_N(AXI_ARESET_N[`getvec(1,19)]),
    .AXI_19_ARADDR(AXI_ARADDR[`getvec(33,19)]),
    .AXI_19_ARBURST(AXI_ARBURST[`getvec(2,19)]),
    .AXI_19_ARID(AXI_ARID[`getvec(6,19)]),
    .AXI_19_ARLEN(AXI_ARLEN[`getvec(4,19)]),
    .AXI_19_ARSIZE(AXI_ARSIZE[`getvec(3,19)]),
    .AXI_19_ARVALID(AXI_ARVALID[`getvec(1,19)]),
    .AXI_19_AWADDR(AXI_AWADDR[`getvec(33,19)]),
    .AXI_19_AWBURST(AXI_AWBURST[`getvec(2,19)]),
    .AXI_19_AWID(AXI_AWID[`getvec(6,19)]),
    .AXI_19_AWLEN(AXI_AWLEN[`getvec(4,19)]),
    .AXI_19_AWSIZE(AXI_AWSIZE[`getvec(3,19)]),
    .AXI_19_AWVALID(AXI_AWVALID[`getvec(1,19)]),
    .AXI_19_RREADY(AXI_RREADY[`getvec(1,19)]),
    .AXI_19_BREADY(AXI_BREADY[`getvec(1,19)]),
    .AXI_19_WDATA(AXI_WDATA[`getvec(256,19)]),
    .AXI_19_WLAST(AXI_WLAST[`getvec(1,19)]),
    .AXI_19_WSTRB(AXI_WSTRB[`getvec(32,19)]),
    .AXI_19_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,19)]),
    .AXI_19_WVALID(AXI_WVALID[`getvec(1,19)]),
    .AXI_19_ARREADY(AXI_ARREADY[`getvec(1,19)]),
    .AXI_19_AWREADY(AXI_AWREADY[`getvec(1,19)]),
    .AXI_19_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,19)]),
    .AXI_19_RDATA(AXI_RDATA[`getvec(256,19)]),
    .AXI_19_RID(AXI_RID[`getvec(6,19)]),
    .AXI_19_RLAST(AXI_RLAST[`getvec(1,19)]),
    .AXI_19_RRESP(AXI_RRESP[`getvec(2,19)]),
    .AXI_19_RVALID(AXI_RVALID[`getvec(1,19)]),
    .AXI_19_WREADY(AXI_WREADY[`getvec(1,19)]),
    .AXI_19_BID(AXI_BID[`getvec(6,19)]),
    .AXI_19_BRESP(AXI_BRESP[`getvec(2,19)]),
    .AXI_19_BVALID(AXI_BVALID[`getvec(1,19)]),
    .AXI_20_ACLK(AXI_ACLK[`getvec(1,20)]),
    .AXI_20_ARESET_N(AXI_ARESET_N[`getvec(1,20)]),
    .AXI_20_ARADDR(AXI_ARADDR[`getvec(33,20)]),
    .AXI_20_ARBURST(AXI_ARBURST[`getvec(2,20)]),
    .AXI_20_ARID(AXI_ARID[`getvec(6,20)]),
    .AXI_20_ARLEN(AXI_ARLEN[`getvec(4,20)]),
    .AXI_20_ARSIZE(AXI_ARSIZE[`getvec(3,20)]),
    .AXI_20_ARVALID(AXI_ARVALID[`getvec(1,20)]),
    .AXI_20_AWADDR(AXI_AWADDR[`getvec(33,20)]),
    .AXI_20_AWBURST(AXI_AWBURST[`getvec(2,20)]),
    .AXI_20_AWID(AXI_AWID[`getvec(6,20)]),
    .AXI_20_AWLEN(AXI_AWLEN[`getvec(4,20)]),
    .AXI_20_AWSIZE(AXI_AWSIZE[`getvec(3,20)]),
    .AXI_20_AWVALID(AXI_AWVALID[`getvec(1,20)]),
    .AXI_20_RREADY(AXI_RREADY[`getvec(1,20)]),
    .AXI_20_BREADY(AXI_BREADY[`getvec(1,20)]),
    .AXI_20_WDATA(AXI_WDATA[`getvec(256,20)]),
    .AXI_20_WLAST(AXI_WLAST[`getvec(1,20)]),
    .AXI_20_WSTRB(AXI_WSTRB[`getvec(32,20)]),
    .AXI_20_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,20)]),
    .AXI_20_WVALID(AXI_WVALID[`getvec(1,20)]),
    .AXI_20_ARREADY(AXI_ARREADY[`getvec(1,20)]),
    .AXI_20_AWREADY(AXI_AWREADY[`getvec(1,20)]),
    .AXI_20_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,20)]),
    .AXI_20_RDATA(AXI_RDATA[`getvec(256,20)]),
    .AXI_20_RID(AXI_RID[`getvec(6,20)]),
    .AXI_20_RLAST(AXI_RLAST[`getvec(1,20)]),
    .AXI_20_RRESP(AXI_RRESP[`getvec(2,20)]),
    .AXI_20_RVALID(AXI_RVALID[`getvec(1,20)]),
    .AXI_20_WREADY(AXI_WREADY[`getvec(1,20)]),
    .AXI_20_BID(AXI_BID[`getvec(6,20)]),
    .AXI_20_BRESP(AXI_BRESP[`getvec(2,20)]),
    .AXI_20_BVALID(AXI_BVALID[`getvec(1,20)]),
    .AXI_21_ACLK(AXI_ACLK[`getvec(1,21)]),
    .AXI_21_ARESET_N(AXI_ARESET_N[`getvec(1,21)]),
    .AXI_21_ARADDR(AXI_ARADDR[`getvec(33,21)]),
    .AXI_21_ARBURST(AXI_ARBURST[`getvec(2,21)]),
    .AXI_21_ARID(AXI_ARID[`getvec(6,21)]),
    .AXI_21_ARLEN(AXI_ARLEN[`getvec(4,21)]),
    .AXI_21_ARSIZE(AXI_ARSIZE[`getvec(3,21)]),
    .AXI_21_ARVALID(AXI_ARVALID[`getvec(1,21)]),
    .AXI_21_AWADDR(AXI_AWADDR[`getvec(33,21)]),
    .AXI_21_AWBURST(AXI_AWBURST[`getvec(2,21)]),
    .AXI_21_AWID(AXI_AWID[`getvec(6,21)]),
    .AXI_21_AWLEN(AXI_AWLEN[`getvec(4,21)]),
    .AXI_21_AWSIZE(AXI_AWSIZE[`getvec(3,21)]),
    .AXI_21_AWVALID(AXI_AWVALID[`getvec(1,21)]),
    .AXI_21_RREADY(AXI_RREADY[`getvec(1,21)]),
    .AXI_21_BREADY(AXI_BREADY[`getvec(1,21)]),
    .AXI_21_WDATA(AXI_WDATA[`getvec(256,21)]),
    .AXI_21_WLAST(AXI_WLAST[`getvec(1,21)]),
    .AXI_21_WSTRB(AXI_WSTRB[`getvec(32,21)]),
    .AXI_21_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,21)]),
    .AXI_21_WVALID(AXI_WVALID[`getvec(1,21)]),
    .AXI_21_ARREADY(AXI_ARREADY[`getvec(1,21)]),
    .AXI_21_AWREADY(AXI_AWREADY[`getvec(1,21)]),
    .AXI_21_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,21)]),
    .AXI_21_RDATA(AXI_RDATA[`getvec(256,21)]),
    .AXI_21_RID(AXI_RID[`getvec(6,21)]),
    .AXI_21_RLAST(AXI_RLAST[`getvec(1,21)]),
    .AXI_21_RRESP(AXI_RRESP[`getvec(2,21)]),
    .AXI_21_RVALID(AXI_RVALID[`getvec(1,21)]),
    .AXI_21_WREADY(AXI_WREADY[`getvec(1,21)]),
    .AXI_21_BID(AXI_BID[`getvec(6,21)]),
    .AXI_21_BRESP(AXI_BRESP[`getvec(2,21)]),
    .AXI_21_BVALID(AXI_BVALID[`getvec(1,21)]),
    .AXI_22_ACLK(AXI_ACLK[`getvec(1,22)]),
    .AXI_22_ARESET_N(AXI_ARESET_N[`getvec(1,22)]),
    .AXI_22_ARADDR(AXI_ARADDR[`getvec(33,22)]),
    .AXI_22_ARBURST(AXI_ARBURST[`getvec(2,22)]),
    .AXI_22_ARID(AXI_ARID[`getvec(6,22)]),
    .AXI_22_ARLEN(AXI_ARLEN[`getvec(4,22)]),
    .AXI_22_ARSIZE(AXI_ARSIZE[`getvec(3,22)]),
    .AXI_22_ARVALID(AXI_ARVALID[`getvec(1,22)]),
    .AXI_22_AWADDR(AXI_AWADDR[`getvec(33,22)]),
    .AXI_22_AWBURST(AXI_AWBURST[`getvec(2,22)]),
    .AXI_22_AWID(AXI_AWID[`getvec(6,22)]),
    .AXI_22_AWLEN(AXI_AWLEN[`getvec(4,22)]),
    .AXI_22_AWSIZE(AXI_AWSIZE[`getvec(3,22)]),
    .AXI_22_AWVALID(AXI_AWVALID[`getvec(1,22)]),
    .AXI_22_RREADY(AXI_RREADY[`getvec(1,22)]),
    .AXI_22_BREADY(AXI_BREADY[`getvec(1,22)]),
    .AXI_22_WDATA(AXI_WDATA[`getvec(256,22)]),
    .AXI_22_WLAST(AXI_WLAST[`getvec(1,22)]),
    .AXI_22_WSTRB(AXI_WSTRB[`getvec(32,22)]),
    .AXI_22_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,22)]),
    .AXI_22_WVALID(AXI_WVALID[`getvec(1,22)]),
    .AXI_22_ARREADY(AXI_ARREADY[`getvec(1,22)]),
    .AXI_22_AWREADY(AXI_AWREADY[`getvec(1,22)]),
    .AXI_22_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,22)]),
    .AXI_22_RDATA(AXI_RDATA[`getvec(256,22)]),
    .AXI_22_RID(AXI_RID[`getvec(6,22)]),
    .AXI_22_RLAST(AXI_RLAST[`getvec(1,22)]),
    .AXI_22_RRESP(AXI_RRESP[`getvec(2,22)]),
    .AXI_22_RVALID(AXI_RVALID[`getvec(1,22)]),
    .AXI_22_WREADY(AXI_WREADY[`getvec(1,22)]),
    .AXI_22_BID(AXI_BID[`getvec(6,22)]),
    .AXI_22_BRESP(AXI_BRESP[`getvec(2,22)]),
    .AXI_22_BVALID(AXI_BVALID[`getvec(1,22)]),
    .AXI_23_ACLK(AXI_ACLK[`getvec(1,23)]),
    .AXI_23_ARESET_N(AXI_ARESET_N[`getvec(1,23)]),
    .AXI_23_ARADDR(AXI_ARADDR[`getvec(33,23)]),
    .AXI_23_ARBURST(AXI_ARBURST[`getvec(2,23)]),
    .AXI_23_ARID(AXI_ARID[`getvec(6,23)]),
    .AXI_23_ARLEN(AXI_ARLEN[`getvec(4,23)]),
    .AXI_23_ARSIZE(AXI_ARSIZE[`getvec(3,23)]),
    .AXI_23_ARVALID(AXI_ARVALID[`getvec(1,23)]),
    .AXI_23_AWADDR(AXI_AWADDR[`getvec(33,23)]),
    .AXI_23_AWBURST(AXI_AWBURST[`getvec(2,23)]),
    .AXI_23_AWID(AXI_AWID[`getvec(6,23)]),
    .AXI_23_AWLEN(AXI_AWLEN[`getvec(4,23)]),
    .AXI_23_AWSIZE(AXI_AWSIZE[`getvec(3,23)]),
    .AXI_23_AWVALID(AXI_AWVALID[`getvec(1,23)]),
    .AXI_23_RREADY(AXI_RREADY[`getvec(1,23)]),
    .AXI_23_BREADY(AXI_BREADY[`getvec(1,23)]),
    .AXI_23_WDATA(AXI_WDATA[`getvec(256,23)]),
    .AXI_23_WLAST(AXI_WLAST[`getvec(1,23)]),
    .AXI_23_WSTRB(AXI_WSTRB[`getvec(32,23)]),
    .AXI_23_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,23)]),
    .AXI_23_WVALID(AXI_WVALID[`getvec(1,23)]),
    .AXI_23_ARREADY(AXI_ARREADY[`getvec(1,23)]),
    .AXI_23_AWREADY(AXI_AWREADY[`getvec(1,23)]),
    .AXI_23_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,23)]),
    .AXI_23_RDATA(AXI_RDATA[`getvec(256,23)]),
    .AXI_23_RID(AXI_RID[`getvec(6,23)]),
    .AXI_23_RLAST(AXI_RLAST[`getvec(1,23)]),
    .AXI_23_RRESP(AXI_RRESP[`getvec(2,23)]),
    .AXI_23_RVALID(AXI_RVALID[`getvec(1,23)]),
    .AXI_23_WREADY(AXI_WREADY[`getvec(1,23)]),
    .AXI_23_BID(AXI_BID[`getvec(6,23)]),
    .AXI_23_BRESP(AXI_BRESP[`getvec(2,23)]),
    .AXI_23_BVALID(AXI_BVALID[`getvec(1,23)]),
    .AXI_24_ACLK(AXI_ACLK[`getvec(1,24)]),
    .AXI_24_ARESET_N(AXI_ARESET_N[`getvec(1,24)]),
    .AXI_24_ARADDR(AXI_ARADDR[`getvec(33,24)]),
    .AXI_24_ARBURST(AXI_ARBURST[`getvec(2,24)]),
    .AXI_24_ARID(AXI_ARID[`getvec(6,24)]),
    .AXI_24_ARLEN(AXI_ARLEN[`getvec(4,24)]),
    .AXI_24_ARSIZE(AXI_ARSIZE[`getvec(3,24)]),
    .AXI_24_ARVALID(AXI_ARVALID[`getvec(1,24)]),
    .AXI_24_AWADDR(AXI_AWADDR[`getvec(33,24)]),
    .AXI_24_AWBURST(AXI_AWBURST[`getvec(2,24)]),
    .AXI_24_AWID(AXI_AWID[`getvec(6,24)]),
    .AXI_24_AWLEN(AXI_AWLEN[`getvec(4,24)]),
    .AXI_24_AWSIZE(AXI_AWSIZE[`getvec(3,24)]),
    .AXI_24_AWVALID(AXI_AWVALID[`getvec(1,24)]),
    .AXI_24_RREADY(AXI_RREADY[`getvec(1,24)]),
    .AXI_24_BREADY(AXI_BREADY[`getvec(1,24)]),
    .AXI_24_WDATA(AXI_WDATA[`getvec(256,24)]),
    .AXI_24_WLAST(AXI_WLAST[`getvec(1,24)]),
    .AXI_24_WSTRB(AXI_WSTRB[`getvec(32,24)]),
    .AXI_24_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,24)]),
    .AXI_24_WVALID(AXI_WVALID[`getvec(1,24)]),
    .AXI_24_ARREADY(AXI_ARREADY[`getvec(1,24)]),
    .AXI_24_AWREADY(AXI_AWREADY[`getvec(1,24)]),
    .AXI_24_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,24)]),
    .AXI_24_RDATA(AXI_RDATA[`getvec(256,24)]),
    .AXI_24_RID(AXI_RID[`getvec(6,24)]),
    .AXI_24_RLAST(AXI_RLAST[`getvec(1,24)]),
    .AXI_24_RRESP(AXI_RRESP[`getvec(2,24)]),
    .AXI_24_RVALID(AXI_RVALID[`getvec(1,24)]),
    .AXI_24_WREADY(AXI_WREADY[`getvec(1,24)]),
    .AXI_24_BID(AXI_BID[`getvec(6,24)]),
    .AXI_24_BRESP(AXI_BRESP[`getvec(2,24)]),
    .AXI_24_BVALID(AXI_BVALID[`getvec(1,24)]),
    .AXI_25_ACLK(AXI_ACLK[`getvec(1,25)]),
    .AXI_25_ARESET_N(AXI_ARESET_N[`getvec(1,25)]),
    .AXI_25_ARADDR(AXI_ARADDR[`getvec(33,25)]),
    .AXI_25_ARBURST(AXI_ARBURST[`getvec(2,25)]),
    .AXI_25_ARID(AXI_ARID[`getvec(6,25)]),
    .AXI_25_ARLEN(AXI_ARLEN[`getvec(4,25)]),
    .AXI_25_ARSIZE(AXI_ARSIZE[`getvec(3,25)]),
    .AXI_25_ARVALID(AXI_ARVALID[`getvec(1,25)]),
    .AXI_25_AWADDR(AXI_AWADDR[`getvec(33,25)]),
    .AXI_25_AWBURST(AXI_AWBURST[`getvec(2,25)]),
    .AXI_25_AWID(AXI_AWID[`getvec(6,25)]),
    .AXI_25_AWLEN(AXI_AWLEN[`getvec(4,25)]),
    .AXI_25_AWSIZE(AXI_AWSIZE[`getvec(3,25)]),
    .AXI_25_AWVALID(AXI_AWVALID[`getvec(1,25)]),
    .AXI_25_RREADY(AXI_RREADY[`getvec(1,25)]),
    .AXI_25_BREADY(AXI_BREADY[`getvec(1,25)]),
    .AXI_25_WDATA(AXI_WDATA[`getvec(256,25)]),
    .AXI_25_WLAST(AXI_WLAST[`getvec(1,25)]),
    .AXI_25_WSTRB(AXI_WSTRB[`getvec(32,25)]),
    .AXI_25_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,25)]),
    .AXI_25_WVALID(AXI_WVALID[`getvec(1,25)]),
    .AXI_25_ARREADY(AXI_ARREADY[`getvec(1,25)]),
    .AXI_25_AWREADY(AXI_AWREADY[`getvec(1,25)]),
    .AXI_25_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,25)]),
    .AXI_25_RDATA(AXI_RDATA[`getvec(256,25)]),
    .AXI_25_RID(AXI_RID[`getvec(6,25)]),
    .AXI_25_RLAST(AXI_RLAST[`getvec(1,25)]),
    .AXI_25_RRESP(AXI_RRESP[`getvec(2,25)]),
    .AXI_25_RVALID(AXI_RVALID[`getvec(1,25)]),
    .AXI_25_WREADY(AXI_WREADY[`getvec(1,25)]),
    .AXI_25_BID(AXI_BID[`getvec(6,25)]),
    .AXI_25_BRESP(AXI_BRESP[`getvec(2,25)]),
    .AXI_25_BVALID(AXI_BVALID[`getvec(1,25)]),
    .AXI_26_ACLK(AXI_ACLK[`getvec(1,26)]),
    .AXI_26_ARESET_N(AXI_ARESET_N[`getvec(1,26)]),
    .AXI_26_ARADDR(AXI_ARADDR[`getvec(33,26)]),
    .AXI_26_ARBURST(AXI_ARBURST[`getvec(2,26)]),
    .AXI_26_ARID(AXI_ARID[`getvec(6,26)]),
    .AXI_26_ARLEN(AXI_ARLEN[`getvec(4,26)]),
    .AXI_26_ARSIZE(AXI_ARSIZE[`getvec(3,26)]),
    .AXI_26_ARVALID(AXI_ARVALID[`getvec(1,26)]),
    .AXI_26_AWADDR(AXI_AWADDR[`getvec(33,26)]),
    .AXI_26_AWBURST(AXI_AWBURST[`getvec(2,26)]),
    .AXI_26_AWID(AXI_AWID[`getvec(6,26)]),
    .AXI_26_AWLEN(AXI_AWLEN[`getvec(4,26)]),
    .AXI_26_AWSIZE(AXI_AWSIZE[`getvec(3,26)]),
    .AXI_26_AWVALID(AXI_AWVALID[`getvec(1,26)]),
    .AXI_26_RREADY(AXI_RREADY[`getvec(1,26)]),
    .AXI_26_BREADY(AXI_BREADY[`getvec(1,26)]),
    .AXI_26_WDATA(AXI_WDATA[`getvec(256,26)]),
    .AXI_26_WLAST(AXI_WLAST[`getvec(1,26)]),
    .AXI_26_WSTRB(AXI_WSTRB[`getvec(32,26)]),
    .AXI_26_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,26)]),
    .AXI_26_WVALID(AXI_WVALID[`getvec(1,26)]),
    .AXI_26_ARREADY(AXI_ARREADY[`getvec(1,26)]),
    .AXI_26_AWREADY(AXI_AWREADY[`getvec(1,26)]),
    .AXI_26_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,26)]),
    .AXI_26_RDATA(AXI_RDATA[`getvec(256,26)]),
    .AXI_26_RID(AXI_RID[`getvec(6,26)]),
    .AXI_26_RLAST(AXI_RLAST[`getvec(1,26)]),
    .AXI_26_RRESP(AXI_RRESP[`getvec(2,26)]),
    .AXI_26_RVALID(AXI_RVALID[`getvec(1,26)]),
    .AXI_26_WREADY(AXI_WREADY[`getvec(1,26)]),
    .AXI_26_BID(AXI_BID[`getvec(6,26)]),
    .AXI_26_BRESP(AXI_BRESP[`getvec(2,26)]),
    .AXI_26_BVALID(AXI_BVALID[`getvec(1,26)]),
    .AXI_27_ACLK(AXI_ACLK[`getvec(1,27)]),
    .AXI_27_ARESET_N(AXI_ARESET_N[`getvec(1,27)]),
    .AXI_27_ARADDR(AXI_ARADDR[`getvec(33,27)]),
    .AXI_27_ARBURST(AXI_ARBURST[`getvec(2,27)]),
    .AXI_27_ARID(AXI_ARID[`getvec(6,27)]),
    .AXI_27_ARLEN(AXI_ARLEN[`getvec(4,27)]),
    .AXI_27_ARSIZE(AXI_ARSIZE[`getvec(3,27)]),
    .AXI_27_ARVALID(AXI_ARVALID[`getvec(1,27)]),
    .AXI_27_AWADDR(AXI_AWADDR[`getvec(33,27)]),
    .AXI_27_AWBURST(AXI_AWBURST[`getvec(2,27)]),
    .AXI_27_AWID(AXI_AWID[`getvec(6,27)]),
    .AXI_27_AWLEN(AXI_AWLEN[`getvec(4,27)]),
    .AXI_27_AWSIZE(AXI_AWSIZE[`getvec(3,27)]),
    .AXI_27_AWVALID(AXI_AWVALID[`getvec(1,27)]),
    .AXI_27_RREADY(AXI_RREADY[`getvec(1,27)]),
    .AXI_27_BREADY(AXI_BREADY[`getvec(1,27)]),
    .AXI_27_WDATA(AXI_WDATA[`getvec(256,27)]),
    .AXI_27_WLAST(AXI_WLAST[`getvec(1,27)]),
    .AXI_27_WSTRB(AXI_WSTRB[`getvec(32,27)]),
    .AXI_27_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,27)]),
    .AXI_27_WVALID(AXI_WVALID[`getvec(1,27)]),
    .AXI_27_ARREADY(AXI_ARREADY[`getvec(1,27)]),
    .AXI_27_AWREADY(AXI_AWREADY[`getvec(1,27)]),
    .AXI_27_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,27)]),
    .AXI_27_RDATA(AXI_RDATA[`getvec(256,27)]),
    .AXI_27_RID(AXI_RID[`getvec(6,27)]),
    .AXI_27_RLAST(AXI_RLAST[`getvec(1,27)]),
    .AXI_27_RRESP(AXI_RRESP[`getvec(2,27)]),
    .AXI_27_RVALID(AXI_RVALID[`getvec(1,27)]),
    .AXI_27_WREADY(AXI_WREADY[`getvec(1,27)]),
    .AXI_27_BID(AXI_BID[`getvec(6,27)]),
    .AXI_27_BRESP(AXI_BRESP[`getvec(2,27)]),
    .AXI_27_BVALID(AXI_BVALID[`getvec(1,27)]),
    .AXI_28_ACLK(AXI_ACLK[`getvec(1,28)]),
    .AXI_28_ARESET_N(AXI_ARESET_N[`getvec(1,28)]),
    .AXI_28_ARADDR(AXI_ARADDR[`getvec(33,28)]),
    .AXI_28_ARBURST(AXI_ARBURST[`getvec(2,28)]),
    .AXI_28_ARID(AXI_ARID[`getvec(6,28)]),
    .AXI_28_ARLEN(AXI_ARLEN[`getvec(4,28)]),
    .AXI_28_ARSIZE(AXI_ARSIZE[`getvec(3,28)]),
    .AXI_28_ARVALID(AXI_ARVALID[`getvec(1,28)]),
    .AXI_28_AWADDR(AXI_AWADDR[`getvec(33,28)]),
    .AXI_28_AWBURST(AXI_AWBURST[`getvec(2,28)]),
    .AXI_28_AWID(AXI_AWID[`getvec(6,28)]),
    .AXI_28_AWLEN(AXI_AWLEN[`getvec(4,28)]),
    .AXI_28_AWSIZE(AXI_AWSIZE[`getvec(3,28)]),
    .AXI_28_AWVALID(AXI_AWVALID[`getvec(1,28)]),
    .AXI_28_RREADY(AXI_RREADY[`getvec(1,28)]),
    .AXI_28_BREADY(AXI_BREADY[`getvec(1,28)]),
    .AXI_28_WDATA(AXI_WDATA[`getvec(256,28)]),
    .AXI_28_WLAST(AXI_WLAST[`getvec(1,28)]),
    .AXI_28_WSTRB(AXI_WSTRB[`getvec(32,28)]),
    .AXI_28_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,28)]),
    .AXI_28_WVALID(AXI_WVALID[`getvec(1,28)]),
    .AXI_28_ARREADY(AXI_ARREADY[`getvec(1,28)]),
    .AXI_28_AWREADY(AXI_AWREADY[`getvec(1,28)]),
    .AXI_28_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,28)]),
    .AXI_28_RDATA(AXI_RDATA[`getvec(256,28)]),
    .AXI_28_RID(AXI_RID[`getvec(6,28)]),
    .AXI_28_RLAST(AXI_RLAST[`getvec(1,28)]),
    .AXI_28_RRESP(AXI_RRESP[`getvec(2,28)]),
    .AXI_28_RVALID(AXI_RVALID[`getvec(1,28)]),
    .AXI_28_WREADY(AXI_WREADY[`getvec(1,28)]),
    .AXI_28_BID(AXI_BID[`getvec(6,28)]),
    .AXI_28_BRESP(AXI_BRESP[`getvec(2,28)]),
    .AXI_28_BVALID(AXI_BVALID[`getvec(1,28)]),
    .AXI_29_ACLK(AXI_ACLK[`getvec(1,29)]),
    .AXI_29_ARESET_N(AXI_ARESET_N[`getvec(1,29)]),
    .AXI_29_ARADDR(AXI_ARADDR[`getvec(33,29)]),
    .AXI_29_ARBURST(AXI_ARBURST[`getvec(2,29)]),
    .AXI_29_ARID(AXI_ARID[`getvec(6,29)]),
    .AXI_29_ARLEN(AXI_ARLEN[`getvec(4,29)]),
    .AXI_29_ARSIZE(AXI_ARSIZE[`getvec(3,29)]),
    .AXI_29_ARVALID(AXI_ARVALID[`getvec(1,29)]),
    .AXI_29_AWADDR(AXI_AWADDR[`getvec(33,29)]),
    .AXI_29_AWBURST(AXI_AWBURST[`getvec(2,29)]),
    .AXI_29_AWID(AXI_AWID[`getvec(6,29)]),
    .AXI_29_AWLEN(AXI_AWLEN[`getvec(4,29)]),
    .AXI_29_AWSIZE(AXI_AWSIZE[`getvec(3,29)]),
    .AXI_29_AWVALID(AXI_AWVALID[`getvec(1,29)]),
    .AXI_29_RREADY(AXI_RREADY[`getvec(1,29)]),
    .AXI_29_BREADY(AXI_BREADY[`getvec(1,29)]),
    .AXI_29_WDATA(AXI_WDATA[`getvec(256,29)]),
    .AXI_29_WLAST(AXI_WLAST[`getvec(1,29)]),
    .AXI_29_WSTRB(AXI_WSTRB[`getvec(32,29)]),
    .AXI_29_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,29)]),
    .AXI_29_WVALID(AXI_WVALID[`getvec(1,29)]),
    .AXI_29_ARREADY(AXI_ARREADY[`getvec(1,29)]),
    .AXI_29_AWREADY(AXI_AWREADY[`getvec(1,29)]),
    .AXI_29_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,29)]),
    .AXI_29_RDATA(AXI_RDATA[`getvec(256,29)]),
    .AXI_29_RID(AXI_RID[`getvec(6,29)]),
    .AXI_29_RLAST(AXI_RLAST[`getvec(1,29)]),
    .AXI_29_RRESP(AXI_RRESP[`getvec(2,29)]),
    .AXI_29_RVALID(AXI_RVALID[`getvec(1,29)]),
    .AXI_29_WREADY(AXI_WREADY[`getvec(1,29)]),
    .AXI_29_BID(AXI_BID[`getvec(6,29)]),
    .AXI_29_BRESP(AXI_BRESP[`getvec(2,29)]),
    .AXI_29_BVALID(AXI_BVALID[`getvec(1,29)]),
    .AXI_30_ACLK(AXI_ACLK[`getvec(1,30)]),
    .AXI_30_ARESET_N(AXI_ARESET_N[`getvec(1,30)]),
    .AXI_30_ARADDR(AXI_ARADDR[`getvec(33,30)]),
    .AXI_30_ARBURST(AXI_ARBURST[`getvec(2,30)]),
    .AXI_30_ARID(AXI_ARID[`getvec(6,30)]),
    .AXI_30_ARLEN(AXI_ARLEN[`getvec(4,30)]),
    .AXI_30_ARSIZE(AXI_ARSIZE[`getvec(3,30)]),
    .AXI_30_ARVALID(AXI_ARVALID[`getvec(1,30)]),
    .AXI_30_AWADDR(AXI_AWADDR[`getvec(33,30)]),
    .AXI_30_AWBURST(AXI_AWBURST[`getvec(2,30)]),
    .AXI_30_AWID(AXI_AWID[`getvec(6,30)]),
    .AXI_30_AWLEN(AXI_AWLEN[`getvec(4,30)]),
    .AXI_30_AWSIZE(AXI_AWSIZE[`getvec(3,30)]),
    .AXI_30_AWVALID(AXI_AWVALID[`getvec(1,30)]),
    .AXI_30_RREADY(AXI_RREADY[`getvec(1,30)]),
    .AXI_30_BREADY(AXI_BREADY[`getvec(1,30)]),
    .AXI_30_WDATA(AXI_WDATA[`getvec(256,30)]),
    .AXI_30_WLAST(AXI_WLAST[`getvec(1,30)]),
    .AXI_30_WSTRB(AXI_WSTRB[`getvec(32,30)]),
    .AXI_30_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,30)]),
    .AXI_30_WVALID(AXI_WVALID[`getvec(1,30)]),
    .AXI_30_ARREADY(AXI_ARREADY[`getvec(1,30)]),
    .AXI_30_AWREADY(AXI_AWREADY[`getvec(1,30)]),
    .AXI_30_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,30)]),
    .AXI_30_RDATA(AXI_RDATA[`getvec(256,30)]),
    .AXI_30_RID(AXI_RID[`getvec(6,30)]),
    .AXI_30_RLAST(AXI_RLAST[`getvec(1,30)]),
    .AXI_30_RRESP(AXI_RRESP[`getvec(2,30)]),
    .AXI_30_RVALID(AXI_RVALID[`getvec(1,30)]),
    .AXI_30_WREADY(AXI_WREADY[`getvec(1,30)]),
    .AXI_30_BID(AXI_BID[`getvec(6,30)]),
    .AXI_30_BRESP(AXI_BRESP[`getvec(2,30)]),
    .AXI_30_BVALID(AXI_BVALID[`getvec(1,30)]),
    .AXI_31_ACLK(AXI_ACLK[`getvec(1,31)]),
    .AXI_31_ARESET_N(AXI_ARESET_N[`getvec(1,31)]),
    .AXI_31_ARADDR(AXI_ARADDR[`getvec(33,31)]),
    .AXI_31_ARBURST(AXI_ARBURST[`getvec(2,31)]),
    .AXI_31_ARID(AXI_ARID[`getvec(6,31)]),
    .AXI_31_ARLEN(AXI_ARLEN[`getvec(4,31)]),
    .AXI_31_ARSIZE(AXI_ARSIZE[`getvec(3,31)]),
    .AXI_31_ARVALID(AXI_ARVALID[`getvec(1,31)]),
    .AXI_31_AWADDR(AXI_AWADDR[`getvec(33,31)]),
    .AXI_31_AWBURST(AXI_AWBURST[`getvec(2,31)]),
    .AXI_31_AWID(AXI_AWID[`getvec(6,31)]),
    .AXI_31_AWLEN(AXI_AWLEN[`getvec(4,31)]),
    .AXI_31_AWSIZE(AXI_AWSIZE[`getvec(3,31)]),
    .AXI_31_AWVALID(AXI_AWVALID[`getvec(1,31)]),
    .AXI_31_RREADY(AXI_RREADY[`getvec(1,31)]),
    .AXI_31_BREADY(AXI_BREADY[`getvec(1,31)]),
    .AXI_31_WDATA(AXI_WDATA[`getvec(256,31)]),
    .AXI_31_WLAST(AXI_WLAST[`getvec(1,31)]),
    .AXI_31_WSTRB(AXI_WSTRB[`getvec(32,31)]),
    .AXI_31_WDATA_PARITY(AXI_WDATA_PARITY[`getvec(32,31)]),
    .AXI_31_WVALID(AXI_WVALID[`getvec(1,31)]),
    .AXI_31_ARREADY(AXI_ARREADY[`getvec(1,31)]),
    .AXI_31_AWREADY(AXI_AWREADY[`getvec(1,31)]),
    .AXI_31_RDATA_PARITY(AXI_RDATA_PARITY[`getvec(32,31)]),
    .AXI_31_RDATA(AXI_RDATA[`getvec(256,31)]),
    .AXI_31_RID(AXI_RID[`getvec(6,31)]),
    .AXI_31_RLAST(AXI_RLAST[`getvec(1,31)]),
    .AXI_31_RRESP(AXI_RRESP[`getvec(2,31)]),
    .AXI_31_RVALID(AXI_RVALID[`getvec(1,31)]),
    .AXI_31_WREADY(AXI_WREADY[`getvec(1,31)]),
    .AXI_31_BID(AXI_BID[`getvec(6,31)]),
    .AXI_31_BRESP(AXI_BRESP[`getvec(2,31)]),
    .AXI_31_BVALID(AXI_BVALID[`getvec(1,31)]),


    .APB_0_PCLK(APB_0_PCLK),                    // input wire APB_0_PCLK
    .APB_0_PRESET_N(APB_0_PRESET_N),            // input wire APB_0_PRESET_N

    .APB_1_PCLK(APB_1_PCLK),                    // input wire APB_1_PCLK
    .APB_1_PRESET_N(APB_1_PRESET_N)            // input wire APB_1_PRESET_N


);


endmodule